// megafunction wizard: %FIR II v17.1%
// GENERATION: XML
// fir.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module fir (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [23:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [21:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_0002 fir_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2022 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="17.1" >
// Retrieval info: 	<generic name="filterType" value="single" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="symmetryMode" value="sym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="50" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="0.04" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone IV E" />
// Retrieval info: 	<generic name="speedGrade" value="medium" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="100000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="24" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="-3.204345703125E-4,6.103515625E-5,-1.678466796875E-4,-7.171630859375E-4,-7.62939453125E-4,-1.983642578125E-4,1.068115234375E-4,-4.425048828125E-4,-0.0011444091796875,-9.002685546875E-4,-1.52587890625E-5,9.1552734375E-5,-0.0010528564453125,-0.0018463134765625,-9.765625E-4,3.204345703125E-4,-1.8310546875E-4,-0.0021514892578125,-0.0026702880859375,-7.171630859375E-4,7.781982421875E-4,-9.765625E-4,-0.0037841796875,-0.0033111572265625,1.068115234375E-4,0.0010986328125,-0.0026092529296875,-0.0058135986328125,-0.003265380859375,0.0015716552734375,8.392333984375E-4,-0.005340576171875,-0.007781982421875,-0.0020294189453125,0.00347900390625,-5.950927734375E-4,-0.0092010498046875,-0.0089874267578125,8.392333984375E-4,0.005340576171875,-0.00390625,-0.0139312744140625,-0.0084686279296875,0.0056915283203125,0.0063323974609375,-0.00994873046875,-0.019073486328125,-0.0048675537109375,0.0128936767578125,0.0051116943359375,-0.020050048828125,-0.023895263671875,0.0042724609375,0.0235748291015625,-9.918212890625E-4,-0.0384674072265625,-0.02764892578125,0.027557373046875,0.0446929931640625,-0.023895263671875,-0.095123291015625,-0.0297088623046875,0.187286376953125,0.388671875,0.388671875,0.187286376953125,-0.0297088623046875,-0.095123291015625,-0.023895263671875,0.0446929931640625,0.027557373046875,-0.02764892578125,-0.0384674072265625,-9.918212890625E-4,0.0235748291015625,0.0042724609375,-0.023895263671875,-0.020050048828125,0.0051116943359375,0.0128936767578125,-0.0048675537109375,-0.019073486328125,-0.00994873046875,0.0063323974609375,0.0056915283203125,-0.0084686279296875,-0.0139312744140625,-0.00390625,0.005340576171875,8.392333984375E-4,-0.0089874267578125,-0.0092010498046875,-5.950927734375E-4,0.00347900390625,-0.0020294189453125,-0.007781982421875,-0.005340576171875,8.392333984375E-4,0.0015716552734375,-0.003265380859375,-0.0058135986328125,-0.0026092529296875,0.0010986328125,1.068115234375E-4,-0.0033111572265625,-0.0037841796875,-9.765625E-4,7.781982421875E-4,-7.171630859375E-4,-0.0026702880859375,-0.0021514892578125,-1.8310546875E-4,3.204345703125E-4,-9.765625E-4,-0.0018463134765625,-0.0010528564453125,9.1552734375E-5,-1.52587890625E-5,-9.002685546875E-4,-0.0011444091796875,-4.425048828125E-4,1.068115234375E-4,-1.983642578125E-4,-7.62939453125E-4,-7.171630859375E-4,-1.678466796875E-4,6.103515625E-5,-3.204345703125E-4" />
// Retrieval info: 	<generic name="coeffSetRealValueImag" value="0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, -0.0530093, -0.04498, 0.0, 0.0749693, 0.159034, 0.224907, 0.249809, 0.224907, 0.159034, 0.0749693, 0.0, -0.04498, -0.0530093, -0.0321283, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="16" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffComplex" value="false" />
// Retrieval info: 	<generic name="karatsuba" value="false" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="trunc" />
// Retrieval info: 	<generic name="outMsbBitRem" value="0" />
// Retrieval info: 	<generic name="outLSBRound" value="trunc" />
// Retrieval info: 	<generic name="outLsbBitRem" value="25" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir.vo
// RELATED_FILES: fir.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, fir_0002_rtl_core.vhd, fir_0002_ast.vhd, fir_0002.vhd
