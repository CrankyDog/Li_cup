library verilog;
use verilog.vl_types.all;
entity i2s_tb is
end i2s_tb;
